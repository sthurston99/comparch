module mux_32to1_64(o, s, i00, i01, i02, i03, i04, i05, i06, i07,
								  i08, i09, i10, i11, i12, i13, i14, i15,
								  i16, i17, i18, i19, i20, i21, i22, i23,
								  i24, i25, i26, i27, i28, i29, i30, i31);
								  
	output reg [63:0] o;
	input [4:0] s;
	input [63:0] i00, i01, i02, i03, i04, i05, i06, i07,
					 i08, i09, i10, i11, i12, i13, i14, i15,
					 i16, i17, i18, i19, i20, i21, i22, i23,
					 i24, i25, i26, i27, i28, i29, i30, i31;
					 
	always @(*) begin
		case(s)
			5'd00 : o <= i00;
			5'd01 : o <= i01;
			5'd02 : o <= i02;
			5'd03 : o <= i03;
			5'd04 : o <= i04;
		   5'd05 : o <= i05;
			5'd06 : o <= i06;
			5'd07 : o <= i07;
			5'd08 : o <= i08;
			5'd09 : o <= i09;
			5'd10 : o <= i10;
			5'd11 : o <= i11;
			5'd12 : o <= i12;
			5'd13 : o <= i13;
			5'd14 : o <= i14;
			5'd15 : o <= i15;
			5'd16 : o <= i16;
			5'd17 : o <= i17;
			5'd18 : o <= i18;
			5'd19 : o <= i19;
			5'd20 : o <= i20;
			5'd21 : o <= i21;
			5'd22 : o <= i22;
			5'd23 : o <= i23;
			5'd24 : o <= i24;
			5'd25 : o <= i25;
			5'd26 : o <= i26;
			5'd27 : o <= i27;
			5'd28 : o <= i28;
			5'd29 : o <= i29;
			5'd30 : o <= i30;
			5'd31 : o <= i31;
		endcase
	end
endmodule
